
.include CMOS_Inv.sub
xM1  vin S vout GND sky130_fd_pr__nfet_01v8 w=.42 l=.5
xM2  vin nS vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5

X1  vdd S nS CMOS_Inv		

Vdd vdd 0 3.3
Vin vin 0 pulse(3.3 0 0s 0s 0s 5us 10us)
Vsel S 0 pulse(0 3.3 0s 0s 0s 10us 20us)

.tran 0.01us 20us

.control
run

plot V(vin)
plot V(S)
plot V(vout)
plot V(nS)

.endc

.end
