* F:\eSim_FOSSEE\switch.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/23/21 17:48:46

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
.lib "sky130_fd_pr\models\sky130.lib.spice" tt

xM1  Net-_M1-Pad1_ digital_input vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
xM5  Net-_M1-Pad1_ digital_input GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5
xM2  Net-_M2-Pad1_ Net-_M1-Pad1_ vdd vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
xM6  Net-_M2-Pad1_ Net-_M1-Pad1_ GND GND sky130_fd_pr__nfet_01v8 w=.42 l=.5
xM3  vout Net-_M1-Pad1_ vin_1 vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
xM7  vout Net-_M1-Pad1_ vin_2 GND sky130_fd_pr__nfet_01v8 w=.42 l=.5
xM4  vin_1 Net-_M2-Pad1_ vout GND sky130_fd_pr__nfet_01v8 w=.42 l=.5
xM8  vin_2 Net-_M2-Pad1_ vout vdd sky130_fd_pr__pfet_01v8 w=1 l=0.5
* U1  vdd digital_input vin_1 vin_2 vout PORT

vdd vdd 0 3.3
vin_1 vin_1 0 2.5
vin_2 vin_2 0 2
vd0 digital_input 0 pulse(0 1.8 0s 0s 0s 5us 10us)

.tran .1us 40us

.control
run
plot V(vout) V(digital_input)

.endc

.end
