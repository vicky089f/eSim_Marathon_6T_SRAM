
.include CMOS_Inv.sub
.include TX_Gate.sub

XI1  VDD Net-_XG1-Pad5_ Net-_XG3-Pad2_ CMOS_Inv		
XI3  VDD Net-_XG3-Pad5_ Q CMOS_Inv		
XI4  VDD Q Net-_XG4-Pad2_ CMOS_Inv		
XI2  VDD Net-_XG3-Pad2_ Net-_XG2-Pad2_ CMOS_Inv		
XG3  VDD Net-_XG3-Pad2_ CLK nCLK Net-_XG3-Pad5_ TX_Gate		
XG4  VDD Net-_XG4-Pad2_ nCLK CLK Net-_XG3-Pad5_ TX_Gate		
XG2  VDD Net-_XG2-Pad2_ CLK nCLK Net-_XG1-Pad5_ TX_Gate		
XG1  VDD D nCLK CLK Net-_XG1-Pad5_ TX_Gate		

VDD VDD 0 3.3
Vclk CLK 0 pulse(0 3.3 5us 0.1us 0.1us 5us 10us)
Vnclk nCLK 0 pulse(3.3 0 5us 0.1us 0.1us 5us 10us)
Vd D 0 pulse(0 3.3 3us 0.1us 0.1us 1us 3us)

.tran 0.01us 30us

.control
run

plot V(CLK) V(nCLK)
plot V(D)
plot V(Q)

.endc
.end
