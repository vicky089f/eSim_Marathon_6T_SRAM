* C:\Users\VIGNESH\eSim-Workspace\SRAM\SRAM.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: 06/24/21 22:04:39

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
.lib "sky130_fd_pr\models\sky130.lib.spice" tt

xM2  VOUT Net-_M1-Pad2_ Net-_M2-Pad3_ Net-_M2-Pad3_ sky130_fd_pr__nfet_01v8 w=.42 l=.5
xM1  VOUT Net-_M1-Pad2_ VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.5
xM4  Net-_M1-Pad2_ VOUT Net-_M2-Pad3_ Net-_M2-Pad3_ sky130_fd_pr__nfet_01v8 w=.42 l=.5
xM3  Net-_M1-Pad2_ VOUT VDD VDD sky130_fd_pr__pfet_01v8 w=1 l=0.5
xM6  BLB WL Net-_M1-Pad2_ GND sky130_fd_pr__nfet_01v8 w=.42 l=.5
xM5  BL WL VOUT GND sky130_fd_pr__nfet_01v8 w=.42 l=.5

VDD VDD 0 3.3
VBL BL 0 pulse(0 3.3 0s 0s 0s 5us 10us)
VBLB BLB 0 pulse(3.3 0 0s 0s 0s 5us 10us)
VWL WL 0 pulse(0 3.3 0s 0s 0s 10us 20us)
* VWL WL 0 3.3


.tran 0.1us 20us

.control
run

plot V(WL) V(VOUT)
.endc

.end
